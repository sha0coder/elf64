module elf64

pub fn load(filename string) {
	
}